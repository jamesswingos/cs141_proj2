module alu
    (
        input logic [31:0] x,
        input logic [31:0] y,
        input logic [2:0] op,
        output logic [31:0] z,
        output logic zero, equal, overflow
    );

    // your code here
endmodule
